magic
tech scmos
magscale 1 2
timestamp 1735751134
<< metal1 >>
rect -66 416 -2 616
rect 840 604 930 616
rect 285 537 300 543
rect 461 537 483 543
rect 189 517 204 523
rect 292 517 323 523
rect 477 523 483 537
rect 829 537 844 543
rect 477 517 515 523
rect 333 497 348 503
rect 541 497 556 503
rect -66 404 24 416
rect -66 16 -2 404
rect 365 317 387 323
rect 381 303 387 317
rect 276 297 323 303
rect 381 297 419 303
rect 564 277 579 283
rect 276 257 291 263
rect 866 216 930 604
rect 840 204 930 216
rect 413 137 428 143
rect 557 137 595 143
rect 397 117 412 123
rect 621 117 636 123
rect 525 97 540 103
rect -66 4 24 16
rect 866 4 930 204
<< m2contact >>
rect 348 616 356 624
rect 204 556 212 564
rect 444 556 452 564
rect 476 556 484 564
rect 556 556 564 564
rect 28 536 36 544
rect 220 536 228 544
rect 236 536 244 544
rect 300 536 308 544
rect 380 536 388 544
rect 412 536 420 544
rect 76 516 84 524
rect 204 516 212 524
rect 268 516 276 524
rect 284 516 292 524
rect 364 516 372 524
rect 396 516 404 524
rect 444 516 452 524
rect 492 536 500 544
rect 540 536 548 544
rect 572 536 580 544
rect 748 536 756 544
rect 780 536 788 544
rect 844 536 852 544
rect 588 516 596 524
rect 700 516 708 524
rect 796 516 804 524
rect 236 496 244 504
rect 348 496 356 504
rect 556 496 564 504
rect 828 496 836 504
rect 76 296 84 304
rect 188 296 196 304
rect 252 296 260 304
rect 268 296 276 304
rect 444 316 452 324
rect 572 316 580 324
rect 460 296 468 304
rect 508 296 516 304
rect 524 296 532 304
rect 604 296 612 304
rect 668 296 676 304
rect 780 296 788 304
rect 28 276 36 284
rect 220 276 228 284
rect 300 276 308 284
rect 396 276 404 284
rect 444 276 452 284
rect 492 276 500 284
rect 540 276 548 284
rect 556 276 564 284
rect 620 276 628 284
rect 652 276 660 284
rect 828 276 836 284
rect 204 256 212 264
rect 268 256 276 264
rect 460 256 468 264
rect 556 256 564 264
rect 636 256 644 264
rect 268 156 276 164
rect 364 156 372 164
rect 540 156 548 164
rect 620 156 628 164
rect 636 156 644 164
rect 28 136 36 144
rect 252 136 260 144
rect 284 136 292 144
rect 300 136 308 144
rect 348 136 356 144
rect 428 136 436 144
rect 652 136 660 144
rect 828 136 836 144
rect 76 116 84 124
rect 188 116 196 124
rect 204 116 212 124
rect 236 116 244 124
rect 332 116 340 124
rect 412 116 420 124
rect 444 116 452 124
rect 492 116 500 124
rect 572 116 580 124
rect 636 116 644 124
rect 668 116 676 124
rect 780 116 788 124
rect 380 96 388 104
rect 460 96 468 104
rect 476 96 484 104
rect 540 96 548 104
rect 508 76 516 84
<< metal2 >>
rect 397 657 403 663
rect 189 577 243 583
rect 29 524 35 536
rect 189 524 195 577
rect 205 524 211 556
rect 237 544 243 577
rect 221 524 227 536
rect 301 524 307 536
rect 29 284 35 516
rect 285 503 291 516
rect 349 504 355 616
rect 413 583 419 596
rect 397 577 419 583
rect 397 563 403 577
rect 445 564 451 596
rect 541 577 579 583
rect 388 557 403 563
rect 413 544 419 556
rect 541 544 547 577
rect 573 563 579 577
rect 573 557 588 563
rect 381 524 387 536
rect 244 497 291 503
rect 365 483 371 516
rect 365 477 380 483
rect 397 463 403 516
rect 381 457 403 463
rect 77 304 83 396
rect 189 304 195 316
rect 221 284 227 316
rect 253 304 259 356
rect 269 304 275 316
rect 269 283 275 296
rect 253 277 275 283
rect 29 144 35 276
rect 205 244 211 256
rect 205 143 211 236
rect 253 144 259 277
rect 269 244 275 256
rect 269 164 275 236
rect 285 144 291 196
rect 301 183 307 276
rect 301 177 323 183
rect 189 137 211 143
rect 189 124 195 137
rect 164 117 179 123
rect 173 103 179 117
rect 205 103 211 116
rect 173 97 211 103
rect 237 84 243 116
rect 237 -23 243 76
rect 301 -17 307 136
rect 317 124 323 177
rect 365 164 371 436
rect 381 204 387 457
rect 413 283 419 536
rect 493 524 499 536
rect 557 524 563 556
rect 429 303 435 436
rect 445 324 451 516
rect 525 483 531 516
rect 557 484 563 496
rect 525 477 547 483
rect 461 304 467 396
rect 429 297 451 303
rect 445 284 451 297
rect 493 284 499 316
rect 509 304 515 396
rect 525 304 531 356
rect 541 284 547 477
rect 557 284 563 396
rect 573 324 579 536
rect 701 524 707 556
rect 605 304 611 356
rect 653 284 659 516
rect 404 277 419 283
rect 605 277 620 283
rect 445 257 460 263
rect 349 123 355 136
rect 340 117 355 123
rect 381 104 387 196
rect 413 124 419 196
rect 429 84 435 136
rect 445 124 451 257
rect 557 164 563 256
rect 605 244 611 277
rect 461 104 467 156
rect 541 123 547 156
rect 605 124 611 236
rect 621 164 627 196
rect 637 183 643 256
rect 669 244 675 296
rect 637 177 659 183
rect 653 164 659 177
rect 660 157 675 163
rect 637 143 643 156
rect 621 137 643 143
rect 525 117 547 123
rect 477 104 483 116
rect 493 84 499 116
rect 509 -17 515 76
rect 525 -17 531 117
rect 621 103 627 137
rect 573 97 627 103
rect 541 84 547 96
rect 573 84 579 97
rect 653 84 659 136
rect 669 124 675 157
rect 685 124 691 476
rect 749 404 755 536
rect 781 524 787 536
rect 797 444 803 516
rect 829 484 835 496
rect 781 304 787 356
rect 829 284 835 396
rect 845 364 851 536
rect 829 144 835 276
rect 781 84 787 116
rect 301 -23 323 -17
rect 509 -23 531 -17
<< m3contact >>
rect 204 556 212 564
rect 28 516 36 524
rect 76 516 84 524
rect 188 516 196 524
rect 220 516 228 524
rect 268 516 276 524
rect 300 516 308 524
rect 412 596 420 604
rect 444 596 452 604
rect 380 556 388 564
rect 412 556 420 564
rect 476 556 484 564
rect 556 556 564 564
rect 588 556 596 564
rect 700 556 708 564
rect 380 516 388 524
rect 380 476 388 484
rect 364 436 372 444
rect 76 396 84 404
rect 252 356 260 364
rect 188 316 196 324
rect 220 316 228 324
rect 268 316 276 324
rect 28 276 36 284
rect 204 236 212 244
rect 268 236 276 244
rect 284 196 292 204
rect 76 116 84 124
rect 156 116 164 124
rect 236 76 244 84
rect 492 516 500 524
rect 524 516 532 524
rect 556 516 564 524
rect 428 436 436 444
rect 460 396 468 404
rect 508 396 516 404
rect 444 316 452 324
rect 492 316 500 324
rect 524 356 532 364
rect 556 476 564 484
rect 556 396 564 404
rect 588 516 596 524
rect 652 516 660 524
rect 604 356 612 364
rect 684 476 692 484
rect 380 196 388 204
rect 412 196 420 204
rect 316 116 324 124
rect 604 236 612 244
rect 460 156 468 164
rect 556 156 564 164
rect 476 116 484 124
rect 620 196 628 204
rect 668 236 676 244
rect 652 156 660 164
rect 428 76 436 84
rect 492 76 500 84
rect 572 116 580 124
rect 604 116 612 124
rect 636 116 644 124
rect 780 516 788 524
rect 828 476 836 484
rect 796 436 804 444
rect 748 396 756 404
rect 828 396 836 404
rect 780 356 788 364
rect 844 356 852 364
rect 828 276 836 284
rect 684 116 692 124
rect 540 76 548 84
rect 572 76 580 84
rect 652 76 660 84
rect 780 76 788 84
<< metal3 >>
rect 410 605 422 606
rect 442 605 454 606
rect 410 604 454 605
rect 410 596 412 604
rect 420 596 444 604
rect 452 596 454 604
rect 410 595 454 596
rect 410 594 422 595
rect 442 594 454 595
rect 202 565 214 566
rect 378 565 390 566
rect 202 564 390 565
rect 202 556 204 564
rect 212 556 380 564
rect 388 556 390 564
rect 202 555 390 556
rect 202 554 214 555
rect 378 554 390 555
rect 410 565 422 566
rect 474 565 486 566
rect 554 565 566 566
rect 410 564 566 565
rect 410 556 412 564
rect 420 556 476 564
rect 484 556 556 564
rect 564 556 566 564
rect 410 555 566 556
rect 410 554 422 555
rect 474 554 486 555
rect 554 554 566 555
rect 586 565 598 566
rect 698 565 710 566
rect 586 564 710 565
rect 586 556 588 564
rect 596 556 700 564
rect 708 556 710 564
rect 586 555 710 556
rect 586 554 598 555
rect 698 554 710 555
rect 26 525 38 526
rect -37 524 38 525
rect -37 516 28 524
rect 36 516 38 524
rect -37 515 38 516
rect -37 495 -27 515
rect 26 514 38 515
rect 74 525 86 526
rect 186 525 198 526
rect 74 524 198 525
rect 74 516 76 524
rect 84 516 188 524
rect 196 516 198 524
rect 74 515 198 516
rect 74 514 86 515
rect 186 514 198 515
rect 218 525 230 526
rect 266 525 278 526
rect 218 524 278 525
rect 218 516 220 524
rect 228 516 268 524
rect 276 516 278 524
rect 218 515 278 516
rect 218 514 230 515
rect 266 514 278 515
rect 298 525 310 526
rect 378 525 390 526
rect 490 525 502 526
rect 522 525 534 526
rect 298 524 534 525
rect 298 516 300 524
rect 308 516 380 524
rect 388 516 492 524
rect 500 516 524 524
rect 532 516 534 524
rect 298 515 534 516
rect 298 514 310 515
rect 378 514 390 515
rect 490 514 502 515
rect 522 514 534 515
rect 554 525 566 526
rect 586 525 598 526
rect 554 524 598 525
rect 554 516 556 524
rect 564 516 588 524
rect 596 516 598 524
rect 554 515 598 516
rect 554 514 566 515
rect 586 514 598 515
rect 650 525 662 526
rect 778 525 790 526
rect 650 524 790 525
rect 650 516 652 524
rect 660 516 780 524
rect 788 516 790 524
rect 650 515 790 516
rect 650 514 662 515
rect 778 514 790 515
rect 378 485 390 486
rect 554 485 566 486
rect 378 484 566 485
rect 378 476 380 484
rect 388 476 556 484
rect 564 476 566 484
rect 378 475 566 476
rect 378 474 390 475
rect 554 474 566 475
rect 682 485 694 486
rect 826 485 838 486
rect 682 484 838 485
rect 682 476 684 484
rect 692 476 828 484
rect 836 476 838 484
rect 682 475 838 476
rect 682 474 694 475
rect 826 474 838 475
rect 362 445 374 446
rect 426 445 438 446
rect 794 445 806 446
rect 362 444 806 445
rect 362 436 364 444
rect 372 436 428 444
rect 436 436 796 444
rect 804 436 806 444
rect 362 435 806 436
rect 362 434 374 435
rect 426 434 438 435
rect 794 434 806 435
rect 74 405 86 406
rect 458 405 470 406
rect 74 404 470 405
rect 74 396 76 404
rect 84 396 460 404
rect 468 396 470 404
rect 74 395 470 396
rect 74 394 86 395
rect 458 394 470 395
rect 506 405 518 406
rect 554 405 566 406
rect 506 404 566 405
rect 506 396 508 404
rect 516 396 556 404
rect 564 396 566 404
rect 506 395 566 396
rect 506 394 518 395
rect 554 394 566 395
rect 746 405 758 406
rect 826 405 838 406
rect 746 404 838 405
rect 746 396 748 404
rect 756 396 828 404
rect 836 396 838 404
rect 746 395 838 396
rect 746 394 758 395
rect 826 394 838 395
rect 250 365 262 366
rect 522 365 534 366
rect 602 365 614 366
rect 250 364 614 365
rect 250 356 252 364
rect 260 356 524 364
rect 532 356 604 364
rect 612 356 614 364
rect 250 355 614 356
rect 250 354 262 355
rect 522 354 534 355
rect 602 354 614 355
rect 778 365 790 366
rect 842 365 854 366
rect 778 364 854 365
rect 778 356 780 364
rect 788 356 844 364
rect 852 356 854 364
rect 778 355 854 356
rect 778 354 790 355
rect 842 354 854 355
rect 186 325 198 326
rect 218 325 230 326
rect 266 325 278 326
rect 186 324 278 325
rect 186 316 188 324
rect 196 316 220 324
rect 228 316 268 324
rect 276 316 278 324
rect 186 315 278 316
rect 186 314 198 315
rect 218 314 230 315
rect 266 314 278 315
rect 442 325 454 326
rect 490 325 502 326
rect 442 324 502 325
rect 442 316 444 324
rect 452 316 492 324
rect 500 316 502 324
rect 442 315 502 316
rect 442 314 454 315
rect 490 314 502 315
rect 26 285 38 286
rect 826 285 838 286
rect 26 284 838 285
rect 26 276 28 284
rect 36 276 828 284
rect 836 276 838 284
rect 26 275 838 276
rect 26 274 38 275
rect 826 274 838 275
rect 202 245 214 246
rect 266 245 278 246
rect 202 244 278 245
rect 202 236 204 244
rect 212 236 268 244
rect 276 236 278 244
rect 202 235 278 236
rect 202 234 214 235
rect 266 234 278 235
rect 602 245 614 246
rect 666 245 678 246
rect 602 244 678 245
rect 602 236 604 244
rect 612 236 668 244
rect 676 236 678 244
rect 602 235 678 236
rect 602 234 614 235
rect 666 234 678 235
rect 282 205 294 206
rect 378 205 390 206
rect 282 204 390 205
rect 282 196 284 204
rect 292 196 380 204
rect 388 196 390 204
rect 282 195 390 196
rect 282 194 294 195
rect 378 194 390 195
rect 410 205 422 206
rect 618 205 630 206
rect 410 204 630 205
rect 410 196 412 204
rect 420 196 620 204
rect 628 196 630 204
rect 410 195 630 196
rect 410 194 422 195
rect 618 194 630 195
rect 458 165 470 166
rect 554 165 566 166
rect 650 165 662 166
rect 458 164 662 165
rect 458 156 460 164
rect 468 156 556 164
rect 564 156 652 164
rect 660 156 662 164
rect 458 155 662 156
rect 458 154 470 155
rect 554 154 566 155
rect 650 154 662 155
rect 74 125 86 126
rect 154 125 166 126
rect 74 124 166 125
rect 74 116 76 124
rect 84 116 156 124
rect 164 116 166 124
rect 74 115 166 116
rect 74 114 86 115
rect 154 114 166 115
rect 314 125 326 126
rect 474 125 486 126
rect 570 125 582 126
rect 602 125 614 126
rect 314 124 614 125
rect 314 116 316 124
rect 324 116 476 124
rect 484 116 572 124
rect 580 116 604 124
rect 612 116 614 124
rect 314 115 614 116
rect 314 114 326 115
rect 474 114 486 115
rect 570 114 582 115
rect 602 114 614 115
rect 634 125 646 126
rect 682 125 694 126
rect 634 124 694 125
rect 634 116 636 124
rect 644 116 684 124
rect 692 116 694 124
rect 634 115 694 116
rect 634 114 646 115
rect 682 114 694 115
rect 234 85 246 86
rect 426 85 438 86
rect 490 85 502 86
rect 234 84 502 85
rect 234 76 236 84
rect 244 76 428 84
rect 436 76 492 84
rect 500 76 502 84
rect 234 75 502 76
rect 234 74 246 75
rect 426 74 438 75
rect 490 74 502 75
rect 538 85 550 86
rect 570 85 582 86
rect 538 84 582 85
rect 538 76 540 84
rect 548 76 572 84
rect 580 76 582 84
rect 538 75 582 76
rect 538 74 550 75
rect 570 74 582 75
rect 650 85 662 86
rect 778 85 790 86
rect 650 84 790 85
rect 650 76 652 84
rect 660 76 780 84
rect 788 76 790 84
rect 650 75 790 76
rect 650 74 662 75
rect 778 74 790 75
use NOR3X1  _23_
timestamp 0
transform 1 0 264 0 1 210
box -4 -6 132 206
use INVX1  _24_
timestamp 0
transform 1 0 264 0 -1 210
box -4 -6 36 206
use AOI21X1  _25_
timestamp 0
transform 1 0 392 0 -1 610
box -4 -6 68 206
use OAI21X1  _26_
timestamp 0
transform 1 0 392 0 1 210
box -4 -6 68 206
use INVX1  _27_
timestamp 0
transform -1 0 376 0 -1 210
box -4 -6 36 206
use INVX1  _28_
timestamp 0
transform 1 0 632 0 1 210
box -4 -6 36 206
use INVX1  _29_
timestamp 0
transform 1 0 536 0 -1 210
box -4 -6 36 206
use NAND2X1  _30_
timestamp 0
transform -1 0 424 0 -1 210
box -4 -6 52 206
use AOI21X1  _31_
timestamp 0
transform 1 0 568 0 -1 210
box -4 -6 68 206
use OAI21X1  _32_
timestamp 0
transform 1 0 776 0 -1 610
box -4 -6 68 206
use OR2X2  _33_
timestamp 0
transform 1 0 200 0 1 210
box -4 -6 68 206
use NOR2X1  _34_
timestamp 0
transform -1 0 568 0 1 210
box -4 -6 52 206
use INVX1  _35_
timestamp 0
transform 1 0 552 0 -1 610
box -4 -6 36 206
use OAI21X1  _36_
timestamp 0
transform -1 0 632 0 1 210
box -4 -6 68 206
use NAND2X1  _37_
timestamp 0
transform 1 0 424 0 -1 210
box -4 -6 52 206
use AOI21X1  _38_
timestamp 0
transform -1 0 520 0 1 210
box -4 -6 68 206
use NAND3X1  _39_
timestamp 0
transform 1 0 472 0 -1 210
box -4 -6 68 206
use INVX1  _40_
timestamp 0
transform 1 0 632 0 -1 210
box -4 -6 36 206
use AND2X2  _41_
timestamp 0
transform -1 0 264 0 -1 210
box -4 -6 68 206
use BUFX2  _42_
timestamp 0
transform -1 0 344 0 -1 210
box -4 -6 52 206
use DFFPOSX1  _43_
timestamp 0
transform -1 0 856 0 1 210
box -4 -6 196 206
use DFFPOSX1  _44_
timestamp 0
transform 1 0 8 0 1 210
box -4 -6 196 206
use DFFPOSX1  _45_
timestamp 0
transform -1 0 856 0 -1 210
box -4 -6 196 206
use DFFPOSX1  _46_
timestamp 0
transform 1 0 8 0 -1 210
box -4 -6 196 206
use INVX1  _47_
timestamp 0
transform -1 0 488 0 -1 610
box -4 -6 36 206
use NAND2X1  _48_
timestamp 0
transform -1 0 392 0 -1 610
box -4 -6 52 206
use OAI21X1  _49_
timestamp 0
transform 1 0 488 0 -1 610
box -4 -6 68 206
use INVX1  _50_
timestamp 0
transform 1 0 200 0 -1 610
box -4 -6 36 206
use NAND2X1  _51_
timestamp 0
transform 1 0 296 0 -1 610
box -4 -6 52 206
use OAI21X1  _52_
timestamp 0
transform -1 0 296 0 -1 610
box -4 -6 68 206
use DFFPOSX1  _53_
timestamp 0
transform -1 0 776 0 -1 610
box -4 -6 196 206
use DFFPOSX1  _54_
timestamp 0
transform 1 0 8 0 -1 610
box -4 -6 196 206
use FILL  FILL12600x6150
timestamp 0
transform -1 0 856 0 -1 610
box -4 -6 20 206
<< labels >>
flabel metal1 s 866 4 930 4 7 FreeSans 16 270 0 0 gnd
port 0 nsew
flabel metal1 s -66 4 -2 4 7 FreeSans 16 270 0 0 vdd
port 1 nsew
flabel metal2 s 397 657 403 663 3 FreeSans 16 90 0 0 DataIn
port 2 nsew
flabel metal2 s 317 -23 323 -17 7 FreeSans 16 270 0 0 Done
port 3 nsew
flabel metal2 s 509 -23 515 -17 7 FreeSans 16 270 0 0 Run
port 4 nsew
flabel metal2 s 237 -23 243 -17 7 FreeSans 16 270 0 0 aResetn
port 5 nsew
flabel metal3 s -37 495 -27 505 7 FreeSans 16 0 0 0 clock
port 6 nsew
<< properties >>
string FIXED_BBOX -48 -40 864 660
<< end >>
