VERSION 5.7 ;
  NOWIREEXTENSIONATPIN ON ;
  DIVIDERCHAR "/" ;
  BUSBITCHARS "[]" ;
MACRO processor_9_bits
  CLASS BLOCK ;
  FOREIGN processor_9_bits ;
  ORIGIN 7.200 6.000 ;
  SIZE 136.800 BY 105.000 ;
  PIN gnd
    USE GROUND ;
    PORT
      LAYER metal1 ;
        RECT 52.200 92.400 53.400 93.600 ;
        RECT 0.600 90.600 139.500 92.400 ;
        RECT 49.800 75.450 51.000 75.600 ;
        RECT 52.200 75.450 53.400 75.600 ;
        RECT 49.800 74.550 53.400 75.450 ;
        RECT 49.800 74.400 51.000 74.550 ;
        RECT 52.200 74.400 53.400 74.550 ;
        RECT 129.900 32.400 139.500 90.600 ;
        RECT 0.600 30.600 139.500 32.400 ;
        RECT 129.900 0.600 139.500 30.600 ;
      LAYER metal2 ;
        RECT 52.200 92.400 53.400 93.600 ;
        RECT 52.350 75.600 53.250 92.400 ;
        RECT 52.200 74.400 53.400 75.600 ;
    END
  END gnd
  PIN vdd
    USE POWER ;
    PORT
      LAYER metal1 ;
        RECT -9.900 62.400 -0.300 92.400 ;
        RECT -9.900 60.600 129.000 62.400 ;
        RECT -9.900 2.400 -0.300 60.600 ;
        RECT -9.900 0.600 129.000 2.400 ;
    END
  END vdd
  PIN DataIn
    PORT
      LAYER metal2 ;
        RECT 59.550 98.550 60.450 99.450 ;
    END
  END DataIn
  PIN Done
    PORT
      LAYER metal1 ;
        RECT 45.000 20.400 46.200 21.600 ;
      LAYER metal2 ;
        RECT 45.000 20.400 46.200 21.600 ;
        RECT 45.150 -2.550 46.050 20.400 ;
        RECT 45.150 -3.450 48.450 -2.550 ;
    END
  END Done
  PIN Run
    PORT
      LAYER metal1 ;
        RECT 81.000 23.400 82.200 24.600 ;
        RECT 76.200 11.400 77.400 12.600 ;
      LAYER metal2 ;
        RECT 81.000 23.400 82.200 24.600 ;
        RECT 81.150 18.450 82.050 23.400 ;
        RECT 78.750 17.550 82.050 18.450 ;
        RECT 76.200 11.400 77.400 12.600 ;
        RECT 76.350 -2.550 77.250 11.400 ;
        RECT 78.750 -2.550 79.650 17.550 ;
        RECT 76.350 -3.450 79.650 -2.550 ;
    END
  END Run
  PIN aResetn
    PORT
      LAYER metal1 ;
        RECT 61.800 21.450 63.000 21.600 ;
        RECT 64.200 21.450 65.400 21.600 ;
        RECT 61.800 20.550 65.400 21.450 ;
        RECT 61.800 20.400 63.000 20.550 ;
        RECT 64.200 20.400 65.400 20.550 ;
        RECT 35.400 17.400 36.600 18.600 ;
        RECT 73.800 17.400 75.000 18.600 ;
      LAYER metal2 ;
        RECT 64.200 20.400 65.400 21.600 ;
        RECT 35.400 17.400 36.600 18.600 ;
        RECT 35.550 12.600 36.450 17.400 ;
        RECT 64.350 12.600 65.250 20.400 ;
        RECT 73.800 17.400 75.000 18.600 ;
        RECT 73.950 12.600 74.850 17.400 ;
        RECT 35.400 11.400 36.600 12.600 ;
        RECT 64.200 11.400 65.400 12.600 ;
        RECT 73.800 11.400 75.000 12.600 ;
        RECT 35.550 -3.450 36.450 11.400 ;
      LAYER metal3 ;
        RECT 35.100 12.750 36.900 12.900 ;
        RECT 63.900 12.750 65.700 12.900 ;
        RECT 73.500 12.750 75.300 12.900 ;
        RECT 35.100 11.250 75.300 12.750 ;
        RECT 35.100 11.100 36.900 11.250 ;
        RECT 63.900 11.100 65.700 11.250 ;
        RECT 73.500 11.100 75.300 11.250 ;
    END
  END aResetn
  PIN clock
    PORT
      LAYER metal1 ;
        RECT 4.200 80.400 5.400 81.600 ;
        RECT 112.200 80.400 113.400 81.600 ;
        RECT 4.200 41.400 5.400 42.600 ;
        RECT 124.200 41.400 125.400 42.600 ;
        RECT 4.200 20.400 5.400 21.600 ;
        RECT 124.200 20.400 125.400 21.600 ;
      LAYER metal2 ;
        RECT 4.200 80.400 5.400 81.600 ;
        RECT 112.200 80.400 113.400 81.600 ;
        RECT 4.350 78.600 5.250 80.400 ;
        RECT 4.200 77.400 5.400 78.600 ;
        RECT 4.350 42.600 5.250 77.400 ;
        RECT 112.350 60.600 113.250 80.400 ;
        RECT 112.200 59.400 113.400 60.600 ;
        RECT 124.200 59.400 125.400 60.600 ;
        RECT 124.350 42.600 125.250 59.400 ;
        RECT 4.200 41.400 5.400 42.600 ;
        RECT 124.200 41.400 125.400 42.600 ;
        RECT 4.350 21.600 5.250 41.400 ;
        RECT 124.350 21.600 125.250 41.400 ;
        RECT 4.200 20.400 5.400 21.600 ;
        RECT 124.200 20.400 125.400 21.600 ;
      LAYER metal3 ;
        RECT 3.900 78.750 5.700 78.900 ;
        RECT -5.550 77.250 5.700 78.750 ;
        RECT -5.550 74.250 -4.050 77.250 ;
        RECT 3.900 77.100 5.700 77.250 ;
        RECT 111.900 60.750 113.700 60.900 ;
        RECT 123.900 60.750 125.700 60.900 ;
        RECT 111.900 59.250 125.700 60.750 ;
        RECT 111.900 59.100 113.700 59.250 ;
        RECT 123.900 59.100 125.700 59.250 ;
        RECT 3.900 42.750 5.700 42.900 ;
        RECT 123.900 42.750 125.700 42.900 ;
        RECT 3.900 41.250 125.700 42.750 ;
        RECT 3.900 41.100 5.700 41.250 ;
        RECT 123.900 41.100 125.700 41.250 ;
    END
  END clock
  OBS
      LAYER metal1 ;
        RECT 1.800 82.500 3.000 89.700 ;
        RECT 4.200 83.700 5.400 89.700 ;
        RECT 8.400 87.600 9.600 89.700 ;
        RECT 6.600 86.700 9.600 87.600 ;
        RECT 12.300 86.700 13.800 89.700 ;
        RECT 15.000 86.700 16.200 89.700 ;
        RECT 17.400 86.700 18.600 89.700 ;
        RECT 21.300 87.600 23.100 89.700 ;
        RECT 21.000 86.700 23.100 87.600 ;
        RECT 6.600 85.500 7.800 86.700 ;
        RECT 15.000 85.800 15.900 86.700 ;
        RECT 9.000 84.600 10.200 85.800 ;
        RECT 11.700 84.900 15.900 85.800 ;
        RECT 21.000 85.500 22.200 86.700 ;
        RECT 11.700 84.600 12.900 84.900 ;
        RECT 3.000 80.400 3.300 81.600 ;
        RECT 9.300 81.300 10.200 84.600 ;
        RECT 25.800 84.000 27.000 89.700 ;
        RECT 23.700 83.100 24.900 83.400 ;
        RECT 28.200 83.100 29.400 89.700 ;
        RECT 30.600 86.700 31.800 89.700 ;
        RECT 30.600 85.500 31.800 85.800 ;
        RECT 30.600 83.400 31.800 84.600 ;
        RECT 23.700 82.200 29.400 83.100 ;
        RECT 33.000 82.500 34.200 89.700 ;
        RECT 35.400 83.700 36.600 89.700 ;
        RECT 37.800 84.000 39.000 89.700 ;
        RECT 40.200 84.900 41.400 89.700 ;
        RECT 42.600 84.000 43.800 89.700 ;
        RECT 37.800 83.700 43.800 84.000 ;
        RECT 45.000 83.700 46.200 89.700 ;
        RECT 48.900 84.600 50.100 89.700 ;
        RECT 47.400 83.700 50.100 84.600 ;
        RECT 53.100 84.600 54.300 89.700 ;
        RECT 53.100 83.700 55.800 84.600 ;
        RECT 57.000 83.700 58.200 89.700 ;
        RECT 60.300 83.700 61.500 89.700 ;
        RECT 64.200 83.700 65.400 89.700 ;
        RECT 66.600 86.700 67.800 89.700 ;
        RECT 66.300 85.500 67.500 85.800 ;
        RECT 35.700 82.500 36.600 83.700 ;
        RECT 38.100 83.100 43.500 83.700 ;
        RECT 45.000 82.500 46.200 82.800 ;
        RECT 17.700 81.300 18.900 81.600 ;
        RECT 6.300 80.400 19.500 81.300 ;
        RECT 7.500 80.100 8.700 80.400 ;
        RECT 5.100 78.600 6.300 78.900 ;
        RECT 5.100 77.700 10.500 78.600 ;
        RECT 11.400 77.400 12.600 78.600 ;
        RECT 1.800 76.500 10.200 76.800 ;
        RECT 1.800 76.200 10.500 76.500 ;
        RECT 1.800 75.900 16.500 76.200 ;
        RECT 1.800 63.300 3.000 75.900 ;
        RECT 9.300 75.300 16.500 75.900 ;
        RECT 4.200 63.300 5.400 75.000 ;
        RECT 6.600 73.500 14.700 74.400 ;
        RECT 6.600 73.200 7.800 73.500 ;
        RECT 13.500 73.200 14.700 73.500 ;
        RECT 15.600 73.500 16.500 75.300 ;
        RECT 18.600 75.600 19.500 80.400 ;
        RECT 28.200 79.500 29.400 82.200 ;
        RECT 33.000 80.400 34.200 81.600 ;
        RECT 35.400 80.400 36.600 81.600 ;
        RECT 37.500 80.400 39.300 81.600 ;
        RECT 41.400 80.700 41.700 82.200 ;
        RECT 42.600 81.450 43.800 81.600 ;
        RECT 45.000 81.450 46.200 81.600 ;
        RECT 42.600 80.550 46.200 81.450 ;
        RECT 42.600 80.400 43.800 80.550 ;
        RECT 45.000 80.400 46.200 80.550 ;
        RECT 21.000 79.200 22.200 79.500 ;
        RECT 21.000 78.300 26.700 79.200 ;
        RECT 25.500 78.000 26.700 78.300 ;
        RECT 28.200 78.450 29.400 78.600 ;
        RECT 30.600 78.450 31.800 78.600 ;
        RECT 28.200 77.550 31.800 78.450 ;
        RECT 28.200 77.400 29.400 77.550 ;
        RECT 30.600 77.400 31.800 77.550 ;
        RECT 23.100 77.100 24.300 77.400 ;
        RECT 23.100 76.500 27.300 77.100 ;
        RECT 23.100 76.200 29.400 76.500 ;
        RECT 18.600 74.700 22.200 75.600 ;
        RECT 17.700 73.500 18.900 73.800 ;
        RECT 15.600 72.600 18.900 73.500 ;
        RECT 21.300 73.200 22.200 74.700 ;
        RECT 21.300 72.000 23.400 73.200 ;
        RECT 11.700 71.100 12.900 71.400 ;
        RECT 15.900 71.100 17.100 71.400 ;
        RECT 6.600 69.300 7.800 70.500 ;
        RECT 11.700 70.200 17.100 71.100 ;
        RECT 15.000 69.300 15.900 70.200 ;
        RECT 21.000 69.300 22.200 70.500 ;
        RECT 6.600 68.400 9.600 69.300 ;
        RECT 8.400 63.300 9.600 68.400 ;
        RECT 12.600 63.300 13.800 69.300 ;
        RECT 15.000 63.300 16.200 69.300 ;
        RECT 17.400 63.300 18.600 69.300 ;
        RECT 21.300 63.300 23.100 69.300 ;
        RECT 25.800 63.300 27.000 75.300 ;
        RECT 28.200 63.300 29.400 76.200 ;
        RECT 30.600 63.300 31.800 69.300 ;
        RECT 33.000 63.300 34.200 79.500 ;
        RECT 35.400 74.400 36.600 75.600 ;
        RECT 38.400 75.300 39.300 80.400 ;
        RECT 40.200 79.500 41.400 79.800 ;
        RECT 47.400 79.500 48.600 83.700 ;
        RECT 54.600 79.500 55.800 83.700 ;
        RECT 57.000 82.500 58.200 82.800 ;
        RECT 57.000 80.400 58.200 81.600 ;
        RECT 61.800 80.400 63.000 81.600 ;
        RECT 61.800 79.200 63.000 79.500 ;
        RECT 40.200 77.400 41.400 78.600 ;
        RECT 42.600 78.450 43.800 78.600 ;
        RECT 47.400 78.450 48.600 78.600 ;
        RECT 42.600 77.550 48.600 78.450 ;
        RECT 42.600 77.400 43.800 77.550 ;
        RECT 47.400 77.400 48.600 77.550 ;
        RECT 54.600 77.400 55.800 78.600 ;
        RECT 59.400 77.400 60.600 78.600 ;
        RECT 64.200 78.300 65.100 83.700 ;
        RECT 66.600 83.400 67.800 84.600 ;
        RECT 69.000 82.500 70.200 89.700 ;
        RECT 71.400 86.700 72.600 89.700 ;
        RECT 71.400 85.500 72.600 85.800 ;
        RECT 71.400 83.400 72.600 84.600 ;
        RECT 73.800 84.000 75.000 89.700 ;
        RECT 76.200 84.900 77.400 89.700 ;
        RECT 78.600 84.000 79.800 89.700 ;
        RECT 73.800 83.700 79.800 84.000 ;
        RECT 81.000 83.700 82.200 89.700 ;
        RECT 83.400 86.700 84.600 89.700 ;
        RECT 83.400 85.500 84.600 85.800 ;
        RECT 74.100 83.100 79.500 83.700 ;
        RECT 81.000 82.500 81.900 83.700 ;
        RECT 83.400 83.400 84.600 84.600 ;
        RECT 85.800 82.500 87.000 89.700 ;
        RECT 88.200 83.100 89.400 89.700 ;
        RECT 90.600 84.000 91.800 89.700 ;
        RECT 94.500 87.600 96.300 89.700 ;
        RECT 94.500 86.700 96.600 87.600 ;
        RECT 99.000 86.700 100.200 89.700 ;
        RECT 101.400 86.700 102.600 89.700 ;
        RECT 103.800 86.700 105.300 89.700 ;
        RECT 108.000 87.600 109.200 89.700 ;
        RECT 108.000 86.700 111.000 87.600 ;
        RECT 95.400 85.500 96.600 86.700 ;
        RECT 101.700 85.800 102.600 86.700 ;
        RECT 101.700 84.900 105.900 85.800 ;
        RECT 104.700 84.600 105.900 84.900 ;
        RECT 107.400 84.600 108.600 85.800 ;
        RECT 109.800 85.500 111.000 86.700 ;
        RECT 92.700 83.100 93.900 83.400 ;
        RECT 88.200 82.200 93.900 83.100 ;
        RECT 69.000 81.450 70.200 81.600 ;
        RECT 69.000 80.550 72.450 81.450 ;
        RECT 69.000 80.400 70.200 80.550 ;
        RECT 61.500 76.800 61.800 78.300 ;
        RECT 64.200 77.400 65.700 78.300 ;
        RECT 66.600 77.400 67.800 78.600 ;
        RECT 38.400 74.400 39.900 75.300 ;
        RECT 36.600 72.600 37.500 73.500 ;
        RECT 36.600 71.400 37.800 72.600 ;
        RECT 36.300 63.300 37.500 69.300 ;
        RECT 38.700 63.300 39.900 74.400 ;
        RECT 42.600 63.300 43.800 75.300 ;
        RECT 45.000 63.300 46.200 69.300 ;
        RECT 47.400 63.300 48.600 76.500 ;
        RECT 49.800 73.200 51.000 73.500 ;
        RECT 52.200 73.200 53.400 73.500 ;
        RECT 49.800 63.300 51.000 69.300 ;
        RECT 52.200 63.300 53.400 69.300 ;
        RECT 54.600 63.300 55.800 76.500 ;
        RECT 66.600 75.300 67.500 76.500 ;
        RECT 59.400 74.400 65.400 75.300 ;
        RECT 57.000 63.300 58.200 69.300 ;
        RECT 59.400 63.300 60.600 74.400 ;
        RECT 61.800 63.300 63.000 73.500 ;
        RECT 64.200 63.300 65.400 74.400 ;
        RECT 66.600 63.300 67.800 75.300 ;
        RECT 69.000 63.300 70.200 79.500 ;
        RECT 71.550 78.450 72.450 80.550 ;
        RECT 73.800 80.400 75.000 81.600 ;
        RECT 75.900 80.700 76.200 82.200 ;
        RECT 78.300 80.400 80.100 81.600 ;
        RECT 81.000 80.400 82.200 81.600 ;
        RECT 85.800 80.400 87.000 81.600 ;
        RECT 76.200 79.500 77.400 79.800 ;
        RECT 76.200 78.450 77.400 78.600 ;
        RECT 71.550 77.550 77.400 78.450 ;
        RECT 76.200 77.400 77.400 77.550 ;
        RECT 78.300 75.300 79.200 80.400 ;
        RECT 88.200 79.500 89.400 82.200 ;
        RECT 98.700 81.300 99.900 81.600 ;
        RECT 107.400 81.300 108.300 84.600 ;
        RECT 112.200 83.700 113.400 89.700 ;
        RECT 114.600 82.500 115.800 89.700 ;
        RECT 117.000 84.000 118.200 89.700 ;
        RECT 119.400 84.900 120.600 89.700 ;
        RECT 121.800 84.000 123.000 89.700 ;
        RECT 117.000 83.700 123.000 84.000 ;
        RECT 124.200 83.700 125.400 89.700 ;
        RECT 117.300 83.100 122.700 83.700 ;
        RECT 124.200 82.500 125.100 83.700 ;
        RECT 98.100 80.400 111.300 81.300 ;
        RECT 114.300 80.400 114.600 81.600 ;
        RECT 117.000 80.400 118.200 81.600 ;
        RECT 119.100 80.700 119.400 82.200 ;
        RECT 121.500 80.400 123.300 81.600 ;
        RECT 124.200 81.450 125.400 81.600 ;
        RECT 126.600 81.450 127.800 81.600 ;
        RECT 124.200 80.550 127.800 81.450 ;
        RECT 124.200 80.400 125.400 80.550 ;
        RECT 126.600 80.400 127.800 80.550 ;
        RECT 71.400 63.300 72.600 69.300 ;
        RECT 73.800 63.300 75.000 75.300 ;
        RECT 77.700 74.400 79.200 75.300 ;
        RECT 81.000 75.450 82.200 75.600 ;
        RECT 83.400 75.450 84.600 75.600 ;
        RECT 81.000 74.550 84.600 75.450 ;
        RECT 81.000 74.400 82.200 74.550 ;
        RECT 83.400 74.400 84.600 74.550 ;
        RECT 77.700 63.300 78.900 74.400 ;
        RECT 80.100 72.600 81.000 73.500 ;
        RECT 79.800 71.400 81.000 72.600 ;
        RECT 80.100 63.300 81.300 69.300 ;
        RECT 83.400 63.300 84.600 69.300 ;
        RECT 85.800 63.300 87.000 79.500 ;
        RECT 95.400 79.200 96.600 79.500 ;
        RECT 88.200 77.400 89.400 78.600 ;
        RECT 90.900 78.300 96.600 79.200 ;
        RECT 90.900 78.000 92.100 78.300 ;
        RECT 93.300 77.100 94.500 77.400 ;
        RECT 90.300 76.500 94.500 77.100 ;
        RECT 88.200 76.200 94.500 76.500 ;
        RECT 88.200 63.300 89.400 76.200 ;
        RECT 98.100 75.600 99.000 80.400 ;
        RECT 108.900 80.100 110.100 80.400 ;
        RECT 119.400 79.500 120.600 79.800 ;
        RECT 111.300 78.600 112.500 78.900 ;
        RECT 105.000 77.400 106.200 78.600 ;
        RECT 107.100 77.700 112.500 78.600 ;
        RECT 119.400 77.400 120.600 78.600 ;
        RECT 107.400 76.500 115.800 76.800 ;
        RECT 107.100 76.200 115.800 76.500 ;
        RECT 90.600 63.300 91.800 75.300 ;
        RECT 95.400 74.700 99.000 75.600 ;
        RECT 101.100 75.900 115.800 76.200 ;
        RECT 101.100 75.300 108.300 75.900 ;
        RECT 95.400 73.200 96.300 74.700 ;
        RECT 94.200 72.000 96.300 73.200 ;
        RECT 98.700 73.500 99.900 73.800 ;
        RECT 101.100 73.500 102.000 75.300 ;
        RECT 98.700 72.600 102.000 73.500 ;
        RECT 102.900 73.500 111.000 74.400 ;
        RECT 102.900 73.200 104.100 73.500 ;
        RECT 109.800 73.200 111.000 73.500 ;
        RECT 100.500 71.100 101.700 71.400 ;
        RECT 104.700 71.100 105.900 71.400 ;
        RECT 95.400 69.300 96.600 70.500 ;
        RECT 100.500 70.200 105.900 71.100 ;
        RECT 101.700 69.300 102.600 70.200 ;
        RECT 109.800 69.300 111.000 70.500 ;
        RECT 94.500 63.300 96.300 69.300 ;
        RECT 99.000 63.300 100.200 69.300 ;
        RECT 101.400 63.300 102.600 69.300 ;
        RECT 103.800 63.300 105.000 69.300 ;
        RECT 108.000 68.400 111.000 69.300 ;
        RECT 108.000 63.300 109.200 68.400 ;
        RECT 112.200 63.300 113.400 75.000 ;
        RECT 114.600 63.300 115.800 75.900 ;
        RECT 121.500 75.300 122.400 80.400 ;
        RECT 117.000 63.300 118.200 75.300 ;
        RECT 120.900 74.400 122.400 75.300 ;
        RECT 124.200 74.400 125.400 75.600 ;
        RECT 120.900 63.300 122.100 74.400 ;
        RECT 123.300 72.600 124.200 73.500 ;
        RECT 123.000 71.400 124.200 72.600 ;
        RECT 123.300 63.300 124.500 69.300 ;
        RECT 1.800 47.100 3.000 59.700 ;
        RECT 4.200 48.000 5.400 59.700 ;
        RECT 8.400 54.600 9.600 59.700 ;
        RECT 6.600 53.700 9.600 54.600 ;
        RECT 12.600 53.700 13.800 59.700 ;
        RECT 15.000 53.700 16.200 59.700 ;
        RECT 17.400 53.700 18.600 59.700 ;
        RECT 21.300 53.700 23.100 59.700 ;
        RECT 6.600 52.500 7.800 53.700 ;
        RECT 15.000 52.800 15.900 53.700 ;
        RECT 11.700 51.900 17.100 52.800 ;
        RECT 21.000 52.500 22.200 53.700 ;
        RECT 11.700 51.600 12.900 51.900 ;
        RECT 15.900 51.600 17.100 51.900 ;
        RECT 6.600 49.500 7.800 49.800 ;
        RECT 13.500 49.500 14.700 49.800 ;
        RECT 6.600 48.600 14.700 49.500 ;
        RECT 15.600 49.500 18.900 50.400 ;
        RECT 15.600 47.700 16.500 49.500 ;
        RECT 17.700 49.200 18.900 49.500 ;
        RECT 21.300 49.800 23.400 51.000 ;
        RECT 21.300 48.300 22.200 49.800 ;
        RECT 9.300 47.100 16.500 47.700 ;
        RECT 1.800 46.800 16.500 47.100 ;
        RECT 18.600 47.400 22.200 48.300 ;
        RECT 25.800 47.700 27.000 59.700 ;
        RECT 1.800 46.500 10.500 46.800 ;
        RECT 1.800 46.200 10.200 46.500 ;
        RECT 5.100 44.400 10.500 45.300 ;
        RECT 11.400 44.400 12.600 45.600 ;
        RECT 5.100 44.100 6.300 44.400 ;
        RECT 7.500 42.600 8.700 42.900 ;
        RECT 18.600 42.600 19.500 47.400 ;
        RECT 28.200 46.800 29.400 59.700 ;
        RECT 23.100 46.500 29.400 46.800 ;
        RECT 30.600 46.800 31.800 59.700 ;
        RECT 34.500 47.700 35.700 59.700 ;
        RECT 36.900 48.600 38.100 59.700 ;
        RECT 40.200 50.700 41.400 59.700 ;
        RECT 42.600 50.700 43.800 59.700 ;
        RECT 45.000 58.800 51.000 59.700 ;
        RECT 45.000 50.700 46.200 58.800 ;
        RECT 47.400 50.700 48.600 57.900 ;
        RECT 49.800 51.000 51.000 58.800 ;
        RECT 52.500 58.800 57.900 59.700 ;
        RECT 52.500 58.500 53.400 58.800 ;
        RECT 40.500 49.800 41.400 50.700 ;
        RECT 45.000 49.800 45.900 50.700 ;
        RECT 40.500 48.900 45.900 49.800 ;
        RECT 47.700 50.100 48.600 50.700 ;
        RECT 52.200 50.100 53.400 58.500 ;
        RECT 57.000 58.500 57.900 58.800 ;
        RECT 47.700 49.500 53.400 50.100 ;
        RECT 54.600 49.500 55.800 57.900 ;
        RECT 57.000 49.500 58.200 58.500 ;
        RECT 47.700 49.200 53.100 49.500 ;
        RECT 36.900 47.700 39.000 48.600 ;
        RECT 54.600 48.450 55.800 48.600 ;
        RECT 23.100 45.900 27.300 46.500 ;
        RECT 30.600 46.200 36.600 46.800 ;
        RECT 38.100 46.500 39.000 47.700 ;
        RECT 50.700 47.400 53.700 48.300 ;
        RECT 54.600 47.550 58.050 48.450 ;
        RECT 59.400 47.700 60.600 59.700 ;
        RECT 63.300 48.600 64.500 59.700 ;
        RECT 65.700 53.700 66.900 59.700 ;
        RECT 65.400 50.400 66.600 51.600 ;
        RECT 65.700 49.500 66.600 50.400 ;
        RECT 63.300 47.700 64.800 48.600 ;
        RECT 54.600 47.400 55.800 47.550 ;
        RECT 30.600 45.900 36.900 46.200 ;
        RECT 23.100 45.600 24.300 45.900 ;
        RECT 25.500 44.700 26.700 45.000 ;
        RECT 21.000 43.800 26.700 44.700 ;
        RECT 28.200 44.400 29.400 45.600 ;
        RECT 35.700 45.000 36.900 45.900 ;
        RECT 21.000 43.500 22.200 43.800 ;
        RECT 33.600 43.500 34.800 43.800 ;
        RECT 3.000 41.400 3.300 42.600 ;
        RECT 6.300 41.700 19.500 42.600 ;
        RECT 1.800 33.300 3.000 40.500 ;
        RECT 4.200 33.300 5.400 39.300 ;
        RECT 9.300 38.400 10.200 41.700 ;
        RECT 17.700 41.400 18.900 41.700 ;
        RECT 28.200 40.800 29.400 43.500 ;
        RECT 33.000 41.400 34.200 42.600 ;
        RECT 23.700 39.900 29.400 40.800 ;
        RECT 36.000 40.500 36.900 45.000 ;
        RECT 37.800 44.400 39.000 45.600 ;
        RECT 40.200 45.450 41.400 45.600 ;
        RECT 47.400 45.450 48.600 45.600 ;
        RECT 40.200 44.550 48.600 45.450 ;
        RECT 40.200 44.400 41.400 44.550 ;
        RECT 47.400 44.400 48.600 44.550 ;
        RECT 49.500 44.400 49.800 45.600 ;
        RECT 23.700 39.600 24.900 39.900 ;
        RECT 6.600 36.300 7.800 37.500 ;
        RECT 9.000 37.200 10.200 38.400 ;
        RECT 11.700 38.100 12.900 38.400 ;
        RECT 11.700 37.200 15.900 38.100 ;
        RECT 15.000 36.300 15.900 37.200 ;
        RECT 21.000 36.300 22.200 37.500 ;
        RECT 6.600 35.400 9.600 36.300 ;
        RECT 8.400 33.300 9.600 35.400 ;
        RECT 12.300 33.300 13.800 36.300 ;
        RECT 15.000 33.300 16.200 36.300 ;
        RECT 17.400 33.300 18.600 36.300 ;
        RECT 21.000 35.400 23.100 36.300 ;
        RECT 21.300 33.300 23.100 35.400 ;
        RECT 25.800 33.300 27.000 39.000 ;
        RECT 28.200 33.300 29.400 39.900 ;
        RECT 33.300 39.600 36.900 40.500 ;
        RECT 30.600 38.400 31.800 39.600 ;
        RECT 30.600 37.200 31.800 37.500 ;
        RECT 33.300 36.300 34.200 39.600 ;
        RECT 38.100 39.300 39.000 43.500 ;
        RECT 45.000 41.400 46.200 42.600 ;
        RECT 47.100 41.400 47.400 42.600 ;
        RECT 30.600 33.300 31.800 36.300 ;
        RECT 33.000 33.300 34.200 36.300 ;
        RECT 35.400 33.300 36.600 38.700 ;
        RECT 37.800 33.300 39.000 39.300 ;
        RECT 40.200 39.450 41.400 39.600 ;
        RECT 42.600 39.450 43.800 39.600 ;
        RECT 40.200 38.550 43.800 39.450 ;
        RECT 40.200 38.400 41.400 38.550 ;
        RECT 42.600 38.400 43.800 38.550 ;
        RECT 44.700 38.400 45.300 39.600 ;
        RECT 50.700 37.500 51.600 47.400 ;
        RECT 57.150 45.450 58.050 47.550 ;
        RECT 61.800 45.450 63.000 45.600 ;
        RECT 57.150 44.550 63.000 45.450 ;
        RECT 61.800 44.400 63.000 44.550 ;
        RECT 61.800 43.200 63.000 43.500 ;
        RECT 63.900 42.600 64.800 47.700 ;
        RECT 66.600 47.400 67.800 48.600 ;
        RECT 69.000 47.700 70.200 59.700 ;
        RECT 71.400 48.600 72.600 59.700 ;
        RECT 73.800 49.500 75.000 59.700 ;
        RECT 76.200 48.600 77.400 59.700 ;
        RECT 71.400 47.700 77.400 48.600 ;
        RECT 79.500 48.900 80.700 59.700 ;
        RECT 79.500 47.700 82.200 48.900 ;
        RECT 83.400 47.700 84.600 59.700 ;
        RECT 86.700 53.700 87.900 59.700 ;
        RECT 87.000 50.400 88.200 51.600 ;
        RECT 87.000 49.500 87.900 50.400 ;
        RECT 89.100 48.600 90.300 59.700 ;
        RECT 69.300 46.500 70.200 47.700 ;
        RECT 78.600 46.500 79.800 46.800 ;
        RECT 69.000 44.400 70.200 45.600 ;
        RECT 71.100 44.700 72.600 45.600 ;
        RECT 75.000 44.700 75.300 46.200 ;
        RECT 59.400 41.400 60.600 42.600 ;
        RECT 61.500 40.800 61.800 42.300 ;
        RECT 63.900 41.400 65.700 42.600 ;
        RECT 66.600 41.400 67.800 42.600 ;
        RECT 59.700 39.300 65.100 39.900 ;
        RECT 66.600 39.300 67.500 40.500 ;
        RECT 45.600 36.600 51.600 37.500 ;
        RECT 45.600 36.300 46.500 36.600 ;
        RECT 42.600 33.300 43.800 36.300 ;
        RECT 45.000 35.400 46.500 36.300 ;
        RECT 49.800 36.300 51.600 36.600 ;
        RECT 59.400 39.000 65.400 39.300 ;
        RECT 45.000 33.300 46.200 35.400 ;
        RECT 47.400 33.300 48.600 35.700 ;
        RECT 49.800 33.300 51.000 36.300 ;
        RECT 59.400 33.300 60.600 39.000 ;
        RECT 61.800 33.300 63.000 38.100 ;
        RECT 64.200 33.300 65.400 39.000 ;
        RECT 66.600 33.300 67.800 39.300 ;
        RECT 69.000 38.400 70.200 39.600 ;
        RECT 71.700 39.300 72.600 44.700 ;
        RECT 76.200 44.400 77.400 45.600 ;
        RECT 78.600 44.400 79.800 45.600 ;
        RECT 73.800 43.500 75.000 43.800 ;
        RECT 81.000 43.500 81.900 47.700 ;
        RECT 85.800 47.400 87.000 48.600 ;
        RECT 88.800 47.700 90.300 48.600 ;
        RECT 93.000 47.700 94.200 59.700 ;
        RECT 95.400 53.700 96.600 59.700 ;
        RECT 88.800 42.600 89.700 47.700 ;
        RECT 90.600 44.400 91.800 45.600 ;
        RECT 97.800 43.500 99.000 59.700 ;
        RECT 100.200 46.800 101.400 59.700 ;
        RECT 102.600 47.700 103.800 59.700 ;
        RECT 106.500 53.700 108.300 59.700 ;
        RECT 111.000 53.700 112.200 59.700 ;
        RECT 113.400 53.700 114.600 59.700 ;
        RECT 115.800 53.700 117.000 59.700 ;
        RECT 120.000 54.600 121.200 59.700 ;
        RECT 120.000 53.700 123.000 54.600 ;
        RECT 107.400 52.500 108.600 53.700 ;
        RECT 113.700 52.800 114.600 53.700 ;
        RECT 112.500 51.900 117.900 52.800 ;
        RECT 121.800 52.500 123.000 53.700 ;
        RECT 112.500 51.600 113.700 51.900 ;
        RECT 116.700 51.600 117.900 51.900 ;
        RECT 106.200 49.800 108.300 51.000 ;
        RECT 107.400 48.300 108.300 49.800 ;
        RECT 110.700 49.500 114.000 50.400 ;
        RECT 110.700 49.200 111.900 49.500 ;
        RECT 107.400 47.400 111.000 48.300 ;
        RECT 100.200 46.500 106.500 46.800 ;
        RECT 102.300 45.900 106.500 46.500 ;
        RECT 105.300 45.600 106.500 45.900 ;
        RECT 100.200 44.400 101.400 45.600 ;
        RECT 102.900 44.700 104.100 45.000 ;
        RECT 102.900 43.800 108.600 44.700 ;
        RECT 107.400 43.500 108.600 43.800 ;
        RECT 90.600 43.200 91.800 43.500 ;
        RECT 73.800 41.400 75.000 42.600 ;
        RECT 81.000 41.400 82.200 42.600 ;
        RECT 83.400 42.450 84.600 42.600 ;
        RECT 85.800 42.450 87.000 42.600 ;
        RECT 83.400 41.550 87.000 42.450 ;
        RECT 83.400 41.400 84.600 41.550 ;
        RECT 85.800 41.400 87.000 41.550 ;
        RECT 87.900 41.400 89.700 42.600 ;
        RECT 91.800 40.800 92.100 42.300 ;
        RECT 93.000 41.400 94.200 42.600 ;
        RECT 97.800 41.400 99.000 42.600 ;
        RECT 100.200 40.800 101.400 43.500 ;
        RECT 110.100 42.600 111.000 47.400 ;
        RECT 113.100 47.700 114.000 49.500 ;
        RECT 114.900 49.500 116.100 49.800 ;
        RECT 121.800 49.500 123.000 49.800 ;
        RECT 114.900 48.600 123.000 49.500 ;
        RECT 124.200 48.000 125.400 59.700 ;
        RECT 113.100 47.100 120.300 47.700 ;
        RECT 126.600 47.100 127.800 59.700 ;
        RECT 113.100 46.800 127.800 47.100 ;
        RECT 119.100 46.500 127.800 46.800 ;
        RECT 119.400 46.200 127.800 46.500 ;
        RECT 117.000 44.400 118.200 45.600 ;
        RECT 119.100 44.400 124.500 45.300 ;
        RECT 123.300 44.100 124.500 44.400 ;
        RECT 120.900 42.600 122.100 42.900 ;
        RECT 110.100 41.700 123.300 42.600 ;
        RECT 110.700 41.400 111.900 41.700 ;
        RECT 69.300 37.200 70.500 37.500 ;
        RECT 69.000 33.300 70.200 36.300 ;
        RECT 71.400 33.300 72.600 39.300 ;
        RECT 75.300 33.300 76.500 39.300 ;
        RECT 81.000 36.300 81.900 40.500 ;
        RECT 83.400 38.400 84.600 39.600 ;
        RECT 86.100 39.300 87.000 40.500 ;
        RECT 88.500 39.300 93.900 39.900 ;
        RECT 83.400 37.200 84.600 37.500 ;
        RECT 78.600 33.300 79.800 36.300 ;
        RECT 81.000 33.300 82.200 36.300 ;
        RECT 83.400 33.300 84.600 36.300 ;
        RECT 85.800 33.300 87.000 39.300 ;
        RECT 88.200 39.000 94.200 39.300 ;
        RECT 88.200 33.300 89.400 39.000 ;
        RECT 90.600 33.300 91.800 38.100 ;
        RECT 93.000 33.300 94.200 39.000 ;
        RECT 95.400 38.400 96.600 39.600 ;
        RECT 95.400 37.200 96.600 37.500 ;
        RECT 95.400 33.300 96.600 36.300 ;
        RECT 97.800 33.300 99.000 40.500 ;
        RECT 100.200 39.900 105.900 40.800 ;
        RECT 100.200 33.300 101.400 39.900 ;
        RECT 104.700 39.600 105.900 39.900 ;
        RECT 102.600 33.300 103.800 39.000 ;
        RECT 119.400 38.400 120.300 41.700 ;
        RECT 126.300 41.400 126.600 42.600 ;
        RECT 116.700 38.100 117.900 38.400 ;
        RECT 107.400 36.300 108.600 37.500 ;
        RECT 113.700 37.200 117.900 38.100 ;
        RECT 119.400 37.200 120.600 38.400 ;
        RECT 113.700 36.300 114.600 37.200 ;
        RECT 121.800 36.300 123.000 37.500 ;
        RECT 106.500 35.400 108.600 36.300 ;
        RECT 106.500 33.300 108.300 35.400 ;
        RECT 111.000 33.300 112.200 36.300 ;
        RECT 113.400 33.300 114.600 36.300 ;
        RECT 115.800 33.300 117.300 36.300 ;
        RECT 120.000 35.400 123.000 36.300 ;
        RECT 120.000 33.300 121.200 35.400 ;
        RECT 124.200 33.300 125.400 39.300 ;
        RECT 126.600 33.300 127.800 40.500 ;
        RECT 1.800 22.500 3.000 29.700 ;
        RECT 4.200 23.700 5.400 29.700 ;
        RECT 8.400 27.600 9.600 29.700 ;
        RECT 6.600 26.700 9.600 27.600 ;
        RECT 12.300 26.700 13.800 29.700 ;
        RECT 15.000 26.700 16.200 29.700 ;
        RECT 17.400 26.700 18.600 29.700 ;
        RECT 21.300 27.600 23.100 29.700 ;
        RECT 21.000 26.700 23.100 27.600 ;
        RECT 6.600 25.500 7.800 26.700 ;
        RECT 15.000 25.800 15.900 26.700 ;
        RECT 9.000 24.600 10.200 25.800 ;
        RECT 11.700 24.900 15.900 25.800 ;
        RECT 21.000 25.500 22.200 26.700 ;
        RECT 11.700 24.600 12.900 24.900 ;
        RECT 3.000 20.400 3.300 21.600 ;
        RECT 9.300 21.300 10.200 24.600 ;
        RECT 25.800 24.000 27.000 29.700 ;
        RECT 23.700 23.100 24.900 23.400 ;
        RECT 28.200 23.100 29.400 29.700 ;
        RECT 31.500 25.200 32.700 29.700 ;
        RECT 23.700 22.200 29.400 23.100 ;
        RECT 17.700 21.300 18.900 21.600 ;
        RECT 6.300 20.400 19.500 21.300 ;
        RECT 7.500 20.100 8.700 20.400 ;
        RECT 5.100 18.600 6.300 18.900 ;
        RECT 5.100 17.700 10.500 18.600 ;
        RECT 11.400 17.400 12.600 18.600 ;
        RECT 1.800 16.500 10.200 16.800 ;
        RECT 1.800 16.200 10.500 16.500 ;
        RECT 1.800 15.900 16.500 16.200 ;
        RECT 1.800 3.300 3.000 15.900 ;
        RECT 9.300 15.300 16.500 15.900 ;
        RECT 4.200 3.300 5.400 15.000 ;
        RECT 6.600 13.500 14.700 14.400 ;
        RECT 6.600 13.200 7.800 13.500 ;
        RECT 13.500 13.200 14.700 13.500 ;
        RECT 15.600 13.500 16.500 15.300 ;
        RECT 18.600 15.600 19.500 20.400 ;
        RECT 28.200 19.500 29.400 22.200 ;
        RECT 30.600 23.700 32.700 25.200 ;
        RECT 33.900 24.000 35.100 29.700 ;
        RECT 37.800 23.700 39.000 29.700 ;
        RECT 40.200 26.700 41.400 29.700 ;
        RECT 40.200 25.500 41.400 25.800 ;
        RECT 30.600 19.500 31.500 23.700 ;
        RECT 37.800 23.400 38.700 23.700 ;
        RECT 40.200 23.400 41.400 24.600 ;
        RECT 36.000 22.800 38.700 23.400 ;
        RECT 32.400 22.500 38.700 22.800 ;
        RECT 42.600 22.500 43.800 29.700 ;
        RECT 45.000 22.500 46.200 29.700 ;
        RECT 47.400 23.700 48.600 29.700 ;
        RECT 49.800 22.800 51.000 29.700 ;
        RECT 32.400 21.900 36.900 22.500 ;
        RECT 47.700 21.900 51.000 22.800 ;
        RECT 52.200 22.500 53.400 29.700 ;
        RECT 54.600 26.700 55.800 29.700 ;
        RECT 54.600 25.500 55.800 25.800 ;
        RECT 57.900 24.600 59.100 29.700 ;
        RECT 54.600 23.400 55.800 24.600 ;
        RECT 57.900 23.700 60.600 24.600 ;
        RECT 61.800 23.700 63.000 29.700 ;
        RECT 64.200 23.700 65.400 29.700 ;
        RECT 68.100 24.600 69.300 29.700 ;
        RECT 66.600 23.700 69.300 24.600 ;
        RECT 32.400 21.600 33.600 21.900 ;
        RECT 21.000 19.200 22.200 19.500 ;
        RECT 21.000 18.300 26.700 19.200 ;
        RECT 25.500 18.000 26.700 18.300 ;
        RECT 28.200 17.400 29.400 18.600 ;
        RECT 30.600 17.400 31.800 18.600 ;
        RECT 23.100 17.100 24.300 17.400 ;
        RECT 23.100 16.500 27.300 17.100 ;
        RECT 32.700 16.500 33.600 21.600 ;
        RECT 34.800 20.700 36.000 21.000 ;
        RECT 34.800 19.800 36.300 20.700 ;
        RECT 37.800 20.400 39.000 21.600 ;
        RECT 42.600 20.400 43.800 21.600 ;
        RECT 35.400 19.500 36.300 19.800 ;
        RECT 37.800 19.200 39.000 19.500 ;
        RECT 23.100 16.200 29.400 16.500 ;
        RECT 18.600 14.700 22.200 15.600 ;
        RECT 17.700 13.500 18.900 13.800 ;
        RECT 15.600 12.600 18.900 13.500 ;
        RECT 21.300 13.200 22.200 14.700 ;
        RECT 21.300 12.000 23.400 13.200 ;
        RECT 11.700 11.100 12.900 11.400 ;
        RECT 15.900 11.100 17.100 11.400 ;
        RECT 6.600 9.300 7.800 10.500 ;
        RECT 11.700 10.200 17.100 11.100 ;
        RECT 15.000 9.300 15.900 10.200 ;
        RECT 21.000 9.300 22.200 10.500 ;
        RECT 6.600 8.400 9.600 9.300 ;
        RECT 8.400 3.300 9.600 8.400 ;
        RECT 12.600 3.300 13.800 9.300 ;
        RECT 15.000 3.300 16.200 9.300 ;
        RECT 17.400 3.300 18.600 9.300 ;
        RECT 21.300 3.300 23.100 9.300 ;
        RECT 25.800 3.300 27.000 15.300 ;
        RECT 28.200 3.300 29.400 16.200 ;
        RECT 30.600 15.300 31.500 16.500 ;
        RECT 32.700 15.600 36.300 16.500 ;
        RECT 30.600 3.300 31.800 15.300 ;
        RECT 33.000 3.300 34.200 14.700 ;
        RECT 35.400 9.300 36.300 15.600 ;
        RECT 35.400 3.300 36.600 9.300 ;
        RECT 37.800 3.300 39.000 9.300 ;
        RECT 40.200 3.300 41.400 9.300 ;
        RECT 42.600 3.300 43.800 19.500 ;
        RECT 45.000 18.600 46.200 19.500 ;
        RECT 45.000 15.300 45.900 18.600 ;
        RECT 47.700 17.400 48.600 21.900 ;
        RECT 52.200 20.400 53.400 21.600 ;
        RECT 49.800 19.500 51.000 19.800 ;
        RECT 59.400 19.500 60.600 23.700 ;
        RECT 61.800 22.500 63.000 22.800 ;
        RECT 64.200 22.500 65.400 22.800 ;
        RECT 66.600 19.500 67.800 23.700 ;
        RECT 71.400 20.700 72.600 29.700 ;
        RECT 76.800 21.300 78.000 29.700 ;
        RECT 81.000 26.700 82.200 29.700 ;
        RECT 81.000 25.500 82.200 25.800 ;
        RECT 83.400 22.500 84.600 29.700 ;
        RECT 86.700 23.700 87.900 29.700 ;
        RECT 90.600 23.700 91.800 29.700 ;
        RECT 93.000 26.700 94.200 29.700 ;
        RECT 95.400 26.700 96.600 29.700 ;
        RECT 92.700 25.500 93.900 25.800 ;
        RECT 95.400 25.500 96.600 25.800 ;
        RECT 83.400 21.450 84.600 21.600 ;
        RECT 88.200 21.450 89.400 21.600 ;
        RECT 76.800 20.700 79.500 21.300 ;
        RECT 77.100 20.400 79.500 20.700 ;
        RECT 83.400 20.550 89.400 21.450 ;
        RECT 83.400 20.400 84.600 20.550 ;
        RECT 88.200 20.400 89.400 20.550 ;
        RECT 49.800 17.400 51.000 18.600 ;
        RECT 46.800 16.200 48.600 17.400 ;
        RECT 47.700 15.300 48.600 16.200 ;
        RECT 45.000 3.300 46.200 15.300 ;
        RECT 47.700 14.400 51.000 15.300 ;
        RECT 47.400 3.300 48.600 13.500 ;
        RECT 49.800 3.300 51.000 14.400 ;
        RECT 52.200 3.300 53.400 19.500 ;
        RECT 59.400 18.450 60.600 18.600 ;
        RECT 61.800 18.450 63.000 18.600 ;
        RECT 59.400 17.550 63.000 18.450 ;
        RECT 59.400 17.400 60.600 17.550 ;
        RECT 61.800 17.400 63.000 17.550 ;
        RECT 66.600 17.400 67.800 18.600 ;
        RECT 75.900 17.400 76.200 18.600 ;
        RECT 71.400 16.500 72.600 16.800 ;
        RECT 78.600 16.500 79.500 20.400 ;
        RECT 57.000 14.400 58.200 15.600 ;
        RECT 57.000 13.200 58.200 13.500 ;
        RECT 54.600 3.300 55.800 9.300 ;
        RECT 57.000 3.300 58.200 9.300 ;
        RECT 59.400 3.300 60.600 16.500 ;
        RECT 61.800 3.300 63.000 9.300 ;
        RECT 64.200 3.300 65.400 9.300 ;
        RECT 66.600 3.300 67.800 16.500 ;
        RECT 69.000 14.400 70.200 15.600 ;
        RECT 71.400 14.400 72.600 15.600 ;
        RECT 78.600 15.450 79.800 15.600 ;
        RECT 81.000 15.450 82.200 15.600 ;
        RECT 78.600 14.550 82.200 15.450 ;
        RECT 78.600 14.400 79.800 14.550 ;
        RECT 81.000 14.400 82.200 14.550 ;
        RECT 76.200 13.500 77.400 13.800 ;
        RECT 69.000 13.200 70.200 13.500 ;
        RECT 78.600 10.500 79.500 13.500 ;
        RECT 74.100 9.600 79.500 10.500 ;
        RECT 74.100 9.300 75.000 9.600 ;
        RECT 69.000 3.300 70.200 9.300 ;
        RECT 71.400 3.300 72.600 9.300 ;
        RECT 73.800 3.300 75.000 9.300 ;
        RECT 78.600 9.300 79.500 9.600 ;
        RECT 76.200 3.300 77.400 8.700 ;
        RECT 78.600 3.300 79.800 9.300 ;
        RECT 81.000 3.300 82.200 9.300 ;
        RECT 83.400 3.300 84.600 19.500 ;
        RECT 88.200 19.200 89.400 19.500 ;
        RECT 85.800 17.400 87.000 18.600 ;
        RECT 90.600 18.300 91.500 23.700 ;
        RECT 93.000 23.400 94.200 24.600 ;
        RECT 95.400 23.400 96.600 24.600 ;
        RECT 97.800 22.500 99.000 29.700 ;
        RECT 100.200 23.100 101.400 29.700 ;
        RECT 102.600 24.000 103.800 29.700 ;
        RECT 106.500 27.600 108.300 29.700 ;
        RECT 106.500 26.700 108.600 27.600 ;
        RECT 111.000 26.700 112.200 29.700 ;
        RECT 113.400 26.700 114.600 29.700 ;
        RECT 115.800 26.700 117.300 29.700 ;
        RECT 120.000 27.600 121.200 29.700 ;
        RECT 120.000 26.700 123.000 27.600 ;
        RECT 107.400 25.500 108.600 26.700 ;
        RECT 113.700 25.800 114.600 26.700 ;
        RECT 113.700 24.900 117.900 25.800 ;
        RECT 116.700 24.600 117.900 24.900 ;
        RECT 119.400 24.600 120.600 25.800 ;
        RECT 121.800 25.500 123.000 26.700 ;
        RECT 104.700 23.100 105.900 23.400 ;
        RECT 100.200 22.200 105.900 23.100 ;
        RECT 97.800 20.400 99.000 21.600 ;
        RECT 100.200 19.500 101.400 22.200 ;
        RECT 110.700 21.300 111.900 21.600 ;
        RECT 119.400 21.300 120.300 24.600 ;
        RECT 124.200 23.700 125.400 29.700 ;
        RECT 126.600 22.500 127.800 29.700 ;
        RECT 110.100 20.400 123.300 21.300 ;
        RECT 126.300 20.400 126.600 21.600 ;
        RECT 93.000 18.450 94.200 18.600 ;
        RECT 95.400 18.450 96.600 18.600 ;
        RECT 87.900 16.800 88.200 18.300 ;
        RECT 90.600 17.400 92.100 18.300 ;
        RECT 93.000 17.550 96.600 18.450 ;
        RECT 93.000 17.400 94.200 17.550 ;
        RECT 95.400 17.400 96.600 17.550 ;
        RECT 93.000 15.300 93.900 16.500 ;
        RECT 85.800 14.400 91.800 15.300 ;
        RECT 85.800 3.300 87.000 14.400 ;
        RECT 88.200 3.300 89.400 13.500 ;
        RECT 90.600 3.300 91.800 14.400 ;
        RECT 93.000 3.300 94.200 15.300 ;
        RECT 95.400 3.300 96.600 9.300 ;
        RECT 97.800 3.300 99.000 19.500 ;
        RECT 107.400 19.200 108.600 19.500 ;
        RECT 100.200 17.400 101.400 18.600 ;
        RECT 102.900 18.300 108.600 19.200 ;
        RECT 102.900 18.000 104.100 18.300 ;
        RECT 105.300 17.100 106.500 17.400 ;
        RECT 102.300 16.500 106.500 17.100 ;
        RECT 100.200 16.200 106.500 16.500 ;
        RECT 100.200 3.300 101.400 16.200 ;
        RECT 110.100 15.600 111.000 20.400 ;
        RECT 120.900 20.100 122.100 20.400 ;
        RECT 123.300 18.600 124.500 18.900 ;
        RECT 117.000 17.400 118.200 18.600 ;
        RECT 119.100 17.700 124.500 18.600 ;
        RECT 119.400 16.500 127.800 16.800 ;
        RECT 119.100 16.200 127.800 16.500 ;
        RECT 102.600 3.300 103.800 15.300 ;
        RECT 107.400 14.700 111.000 15.600 ;
        RECT 113.100 15.900 127.800 16.200 ;
        RECT 113.100 15.300 120.300 15.900 ;
        RECT 107.400 13.200 108.300 14.700 ;
        RECT 106.200 12.000 108.300 13.200 ;
        RECT 110.700 13.500 111.900 13.800 ;
        RECT 113.100 13.500 114.000 15.300 ;
        RECT 110.700 12.600 114.000 13.500 ;
        RECT 114.900 13.500 123.000 14.400 ;
        RECT 114.900 13.200 116.100 13.500 ;
        RECT 121.800 13.200 123.000 13.500 ;
        RECT 112.500 11.100 113.700 11.400 ;
        RECT 116.700 11.100 117.900 11.400 ;
        RECT 107.400 9.300 108.600 10.500 ;
        RECT 112.500 10.200 117.900 11.100 ;
        RECT 113.700 9.300 114.600 10.200 ;
        RECT 121.800 9.300 123.000 10.500 ;
        RECT 106.500 3.300 108.300 9.300 ;
        RECT 111.000 3.300 112.200 9.300 ;
        RECT 113.400 3.300 114.600 9.300 ;
        RECT 115.800 3.300 117.000 9.300 ;
        RECT 120.000 8.400 123.000 9.300 ;
        RECT 120.000 3.300 121.200 8.400 ;
        RECT 124.200 3.300 125.400 15.000 ;
        RECT 126.600 3.300 127.800 15.900 ;
      LAYER metal2 ;
        RECT 61.800 89.400 63.000 90.600 ;
        RECT 66.600 89.400 67.800 90.600 ;
        RECT 61.950 87.450 62.850 89.400 ;
        RECT 1.800 75.300 3.000 83.700 ;
        RECT 6.600 69.300 7.800 86.700 ;
        RECT 11.400 77.400 12.600 78.600 ;
        RECT 21.000 69.300 22.200 86.700 ;
        RECT 28.350 86.550 36.450 87.450 ;
        RECT 28.350 78.600 29.250 86.550 ;
        RECT 30.600 83.400 31.800 84.600 ;
        RECT 30.750 78.600 31.650 83.400 ;
        RECT 35.550 81.600 36.450 86.550 ;
        RECT 59.550 86.550 62.850 87.450 ;
        RECT 57.000 84.450 58.200 84.600 ;
        RECT 59.550 84.450 60.450 86.550 ;
        RECT 66.750 84.600 67.650 89.400 ;
        RECT 81.150 86.550 86.850 87.450 ;
        RECT 57.000 83.550 60.450 84.450 ;
        RECT 57.000 83.400 58.200 83.550 ;
        RECT 61.800 83.400 63.000 84.600 ;
        RECT 66.600 83.400 67.800 84.600 ;
        RECT 71.400 83.400 72.600 84.600 ;
        RECT 61.950 81.600 62.850 83.400 ;
        RECT 81.150 81.600 82.050 86.550 ;
        RECT 83.400 83.400 84.600 84.600 ;
        RECT 85.950 84.450 86.850 86.550 ;
        RECT 88.200 84.450 89.400 84.600 ;
        RECT 85.950 83.550 89.400 84.450 ;
        RECT 88.200 83.400 89.400 83.550 ;
        RECT 33.000 80.400 34.200 81.600 ;
        RECT 35.400 80.400 36.600 81.600 ;
        RECT 45.000 80.400 46.200 81.600 ;
        RECT 57.000 80.400 58.200 81.600 ;
        RECT 61.800 80.400 63.000 81.600 ;
        RECT 73.800 80.400 75.000 81.600 ;
        RECT 81.000 80.400 82.200 81.600 ;
        RECT 33.150 78.600 34.050 80.400 ;
        RECT 45.150 78.600 46.050 80.400 ;
        RECT 57.150 78.600 58.050 80.400 ;
        RECT 28.200 77.400 29.400 78.600 ;
        RECT 30.600 77.400 31.800 78.600 ;
        RECT 33.000 77.400 34.200 78.600 ;
        RECT 40.200 77.400 41.400 78.600 ;
        RECT 42.600 77.400 43.800 78.600 ;
        RECT 45.000 77.400 46.200 78.600 ;
        RECT 54.600 77.400 55.800 78.600 ;
        RECT 57.000 77.400 58.200 78.600 ;
        RECT 59.400 77.400 60.600 78.600 ;
        RECT 35.400 75.450 36.600 75.600 ;
        RECT 42.750 75.450 43.650 77.400 ;
        RECT 35.400 74.550 43.650 75.450 ;
        RECT 35.400 74.400 36.600 74.550 ;
        RECT 54.750 72.450 55.650 77.400 ;
        RECT 57.000 72.450 58.200 72.600 ;
        RECT 54.750 71.550 58.200 72.450 ;
        RECT 57.000 71.400 58.200 71.550 ;
        RECT 59.550 69.450 60.450 77.400 ;
        RECT 57.150 68.550 60.450 69.450 ;
        RECT 54.600 65.400 55.800 66.600 ;
        RECT 11.400 59.400 12.600 60.600 ;
        RECT 1.800 39.300 3.000 47.700 ;
        RECT 6.600 36.300 7.800 53.700 ;
        RECT 11.550 45.600 12.450 59.400 ;
        RECT 11.400 44.400 12.600 45.600 ;
        RECT 21.000 36.300 22.200 53.700 ;
        RECT 37.800 53.400 39.000 54.600 ;
        RECT 28.200 47.400 29.400 48.600 ;
        RECT 33.000 47.400 34.200 48.600 ;
        RECT 28.350 45.600 29.250 47.400 ;
        RECT 28.200 44.400 29.400 45.600 ;
        RECT 33.150 42.600 34.050 47.400 ;
        RECT 37.950 45.600 38.850 53.400 ;
        RECT 40.200 47.400 41.400 48.600 ;
        RECT 40.350 45.600 41.250 47.400 ;
        RECT 37.800 44.400 39.000 45.600 ;
        RECT 40.200 44.400 41.400 45.600 ;
        RECT 33.000 41.400 34.200 42.600 ;
        RECT 40.350 42.450 41.250 44.400 ;
        RECT 37.950 41.550 41.250 42.450 ;
        RECT 30.600 38.400 31.800 39.600 ;
        RECT 30.750 36.600 31.650 38.400 ;
        RECT 30.600 35.400 31.800 36.600 ;
        RECT 1.800 15.300 3.000 23.700 ;
        RECT 6.600 9.300 7.800 26.700 ;
        RECT 11.400 17.400 12.600 18.600 ;
        RECT 21.000 9.300 22.200 26.700 ;
        RECT 30.750 21.450 31.650 35.400 ;
        RECT 37.950 21.600 38.850 41.550 ;
        RECT 45.000 41.400 46.200 42.600 ;
        RECT 40.200 38.400 41.400 39.600 ;
        RECT 40.350 36.600 41.250 38.400 ;
        RECT 40.200 35.400 41.400 36.600 ;
        RECT 40.350 24.600 41.250 35.400 ;
        RECT 42.600 29.400 43.800 30.600 ;
        RECT 40.200 23.400 41.400 24.600 ;
        RECT 42.750 21.600 43.650 29.400 ;
        RECT 45.150 27.450 46.050 41.400 ;
        RECT 45.150 26.550 48.450 27.450 ;
        RECT 28.350 20.550 31.650 21.450 ;
        RECT 28.350 18.600 29.250 20.550 ;
        RECT 37.800 20.400 39.000 21.600 ;
        RECT 42.600 20.400 43.800 21.600 ;
        RECT 47.550 18.600 48.450 26.550 ;
        RECT 54.750 24.600 55.650 65.400 ;
        RECT 57.150 30.600 58.050 68.550 ;
        RECT 59.400 42.450 60.600 42.600 ;
        RECT 61.950 42.450 62.850 80.400 ;
        RECT 73.950 78.600 74.850 80.400 ;
        RECT 83.550 78.600 84.450 83.400 ;
        RECT 85.800 80.400 87.000 81.600 ;
        RECT 66.600 77.400 67.800 78.600 ;
        RECT 73.800 77.400 75.000 78.600 ;
        RECT 78.600 77.400 79.800 78.600 ;
        RECT 83.400 77.400 84.600 78.600 ;
        RECT 64.200 65.400 65.400 66.600 ;
        RECT 64.350 45.450 65.250 65.400 ;
        RECT 66.750 48.600 67.650 77.400 ;
        RECT 78.750 72.450 79.650 77.400 ;
        RECT 83.400 74.400 84.600 75.600 ;
        RECT 83.550 72.600 84.450 74.400 ;
        RECT 78.750 71.550 82.050 72.450 ;
        RECT 69.000 59.400 70.200 60.600 ;
        RECT 76.200 59.400 77.400 60.600 ;
        RECT 66.600 47.400 67.800 48.600 ;
        RECT 69.150 45.600 70.050 59.400 ;
        RECT 73.800 47.400 75.000 48.600 ;
        RECT 64.350 44.550 67.650 45.450 ;
        RECT 66.750 42.600 67.650 44.550 ;
        RECT 69.000 44.400 70.200 45.600 ;
        RECT 73.950 42.600 74.850 47.400 ;
        RECT 76.350 45.600 77.250 59.400 ;
        RECT 78.600 53.400 79.800 54.600 ;
        RECT 78.750 45.600 79.650 53.400 ;
        RECT 76.200 44.400 77.400 45.600 ;
        RECT 78.600 44.400 79.800 45.600 ;
        RECT 81.150 42.600 82.050 71.550 ;
        RECT 83.400 71.400 84.600 72.600 ;
        RECT 83.400 59.400 84.600 60.600 ;
        RECT 83.550 42.600 84.450 59.400 ;
        RECT 85.950 48.600 86.850 80.400 ;
        RECT 88.200 77.400 89.400 78.600 ;
        RECT 95.400 69.300 96.600 86.700 ;
        RECT 105.000 83.400 106.200 84.600 ;
        RECT 105.150 78.600 106.050 83.400 ;
        RECT 97.800 77.400 99.000 78.600 ;
        RECT 105.000 77.400 106.200 78.600 ;
        RECT 90.600 53.400 91.800 54.600 ;
        RECT 85.800 47.400 87.000 48.600 ;
        RECT 90.750 45.600 91.650 53.400 ;
        RECT 90.600 44.400 91.800 45.600 ;
        RECT 97.950 42.600 98.850 77.400 ;
        RECT 102.600 71.400 103.800 72.600 ;
        RECT 100.200 44.400 101.400 45.600 ;
        RECT 59.400 41.550 62.850 42.450 ;
        RECT 59.400 41.400 60.600 41.550 ;
        RECT 66.600 41.400 67.800 42.600 ;
        RECT 73.800 41.400 75.000 42.600 ;
        RECT 81.000 41.400 82.200 42.600 ;
        RECT 83.400 41.400 84.600 42.600 ;
        RECT 93.000 42.450 94.200 42.600 ;
        RECT 90.750 41.550 94.200 42.450 ;
        RECT 69.000 39.450 70.200 39.600 ;
        RECT 66.750 38.550 70.200 39.450 ;
        RECT 57.000 29.400 58.200 30.600 ;
        RECT 61.800 29.400 63.000 30.600 ;
        RECT 54.600 23.400 55.800 24.600 ;
        RECT 52.200 20.400 53.400 21.600 ;
        RECT 23.400 18.450 24.600 18.600 ;
        RECT 23.400 17.550 26.850 18.450 ;
        RECT 23.400 17.400 24.600 17.550 ;
        RECT 25.950 15.450 26.850 17.550 ;
        RECT 28.200 17.400 29.400 18.600 ;
        RECT 30.600 17.400 31.800 18.600 ;
        RECT 47.400 17.400 48.600 18.600 ;
        RECT 49.800 18.450 51.000 18.600 ;
        RECT 52.350 18.450 53.250 20.400 ;
        RECT 49.800 17.550 53.250 18.450 ;
        RECT 49.800 17.400 51.000 17.550 ;
        RECT 30.750 15.450 31.650 17.400 ;
        RECT 57.150 15.600 58.050 29.400 ;
        RECT 61.950 18.600 62.850 29.400 ;
        RECT 66.750 18.600 67.650 38.550 ;
        RECT 69.000 38.400 70.200 38.550 ;
        RECT 83.400 38.400 84.600 39.600 ;
        RECT 83.550 24.600 84.450 38.400 ;
        RECT 90.750 36.600 91.650 41.550 ;
        RECT 93.000 41.400 94.200 41.550 ;
        RECT 97.800 41.400 99.000 42.600 ;
        RECT 95.400 38.400 96.600 39.600 ;
        RECT 90.600 35.400 91.800 36.600 ;
        RECT 69.000 23.400 70.200 24.600 ;
        RECT 83.400 23.400 84.600 24.600 ;
        RECT 61.800 17.400 63.000 18.600 ;
        RECT 66.600 17.400 67.800 18.600 ;
        RECT 69.150 15.600 70.050 23.400 ;
        RECT 90.750 18.600 91.650 35.400 ;
        RECT 93.000 29.400 94.200 30.600 ;
        RECT 93.150 24.600 94.050 29.400 ;
        RECT 95.550 27.450 96.450 38.400 ;
        RECT 100.350 36.600 101.250 44.400 ;
        RECT 100.200 35.400 101.400 36.600 ;
        RECT 95.550 26.550 98.850 27.450 ;
        RECT 97.950 24.600 98.850 26.550 ;
        RECT 93.000 23.400 94.200 24.600 ;
        RECT 95.400 23.400 96.600 24.600 ;
        RECT 97.800 24.450 99.000 24.600 ;
        RECT 97.800 23.550 101.250 24.450 ;
        RECT 97.800 23.400 99.000 23.550 ;
        RECT 95.550 21.450 96.450 23.400 ;
        RECT 93.150 20.550 96.450 21.450 ;
        RECT 71.400 17.400 72.600 18.600 ;
        RECT 85.800 17.400 87.000 18.600 ;
        RECT 90.600 17.400 91.800 18.600 ;
        RECT 71.550 15.600 72.450 17.400 ;
        RECT 25.950 14.550 31.650 15.450 ;
        RECT 57.000 14.400 58.200 15.600 ;
        RECT 69.000 14.400 70.200 15.600 ;
        RECT 71.400 14.400 72.600 15.600 ;
        RECT 81.000 14.400 82.200 15.600 ;
        RECT 93.150 15.450 94.050 20.550 ;
        RECT 97.800 20.400 99.000 21.600 ;
        RECT 95.400 17.400 96.600 18.600 ;
        RECT 85.950 14.550 94.050 15.450 ;
        RECT 81.150 12.600 82.050 14.400 ;
        RECT 85.950 12.600 86.850 14.550 ;
        RECT 97.950 12.600 98.850 20.400 ;
        RECT 100.350 18.600 101.250 23.550 ;
        RECT 102.750 18.600 103.650 71.400 ;
        RECT 109.800 69.300 111.000 86.700 ;
        RECT 114.600 75.300 115.800 83.700 ;
        RECT 117.000 80.400 118.200 81.600 ;
        RECT 126.600 80.400 127.800 81.600 ;
        RECT 117.150 78.600 118.050 80.400 ;
        RECT 117.000 77.400 118.200 78.600 ;
        RECT 119.400 77.400 120.600 78.600 ;
        RECT 119.550 66.600 120.450 77.400 ;
        RECT 124.200 74.400 125.400 75.600 ;
        RECT 124.350 72.600 125.250 74.400 ;
        RECT 124.200 71.400 125.400 72.600 ;
        RECT 119.400 65.400 120.600 66.600 ;
        RECT 126.750 54.600 127.650 80.400 ;
        RECT 107.400 36.300 108.600 53.700 ;
        RECT 117.000 53.400 118.200 54.600 ;
        RECT 117.150 45.600 118.050 53.400 ;
        RECT 117.000 44.400 118.200 45.600 ;
        RECT 121.800 36.300 123.000 53.700 ;
        RECT 126.600 53.400 127.800 54.600 ;
        RECT 126.600 39.300 127.800 47.700 ;
        RECT 100.200 17.400 101.400 18.600 ;
        RECT 102.600 17.400 103.800 18.600 ;
        RECT 81.000 11.400 82.200 12.600 ;
        RECT 85.800 11.400 87.000 12.600 ;
        RECT 97.800 11.400 99.000 12.600 ;
        RECT 107.400 9.300 108.600 26.700 ;
        RECT 117.000 17.400 118.200 18.600 ;
        RECT 117.150 12.600 118.050 17.400 ;
        RECT 117.000 11.400 118.200 12.600 ;
        RECT 121.800 9.300 123.000 26.700 ;
        RECT 126.600 15.300 127.800 23.700 ;
      LAYER metal3 ;
        RECT 61.500 90.750 63.300 90.900 ;
        RECT 66.300 90.750 68.100 90.900 ;
        RECT 61.500 89.250 68.100 90.750 ;
        RECT 61.500 89.100 63.300 89.250 ;
        RECT 66.300 89.100 68.100 89.250 ;
        RECT 30.300 84.750 32.100 84.900 ;
        RECT 56.700 84.750 58.500 84.900 ;
        RECT 30.300 83.250 58.500 84.750 ;
        RECT 30.300 83.100 32.100 83.250 ;
        RECT 56.700 83.100 58.500 83.250 ;
        RECT 61.500 84.750 63.300 84.900 ;
        RECT 71.100 84.750 72.900 84.900 ;
        RECT 83.100 84.750 84.900 84.900 ;
        RECT 61.500 83.250 84.900 84.750 ;
        RECT 61.500 83.100 63.300 83.250 ;
        RECT 71.100 83.100 72.900 83.250 ;
        RECT 83.100 83.100 84.900 83.250 ;
        RECT 87.900 84.750 89.700 84.900 ;
        RECT 104.700 84.750 106.500 84.900 ;
        RECT 87.900 83.250 106.500 84.750 ;
        RECT 87.900 83.100 89.700 83.250 ;
        RECT 104.700 83.100 106.500 83.250 ;
        RECT 11.100 78.750 12.900 78.900 ;
        RECT 27.900 78.750 29.700 78.900 ;
        RECT 11.100 77.250 29.700 78.750 ;
        RECT 11.100 77.100 12.900 77.250 ;
        RECT 27.900 77.100 29.700 77.250 ;
        RECT 32.700 78.750 34.500 78.900 ;
        RECT 39.900 78.750 41.700 78.900 ;
        RECT 32.700 77.250 41.700 78.750 ;
        RECT 32.700 77.100 34.500 77.250 ;
        RECT 39.900 77.100 41.700 77.250 ;
        RECT 44.700 78.750 46.500 78.900 ;
        RECT 56.700 78.750 58.500 78.900 ;
        RECT 73.500 78.750 75.300 78.900 ;
        RECT 78.300 78.750 80.100 78.900 ;
        RECT 44.700 77.250 80.100 78.750 ;
        RECT 44.700 77.100 46.500 77.250 ;
        RECT 56.700 77.100 58.500 77.250 ;
        RECT 73.500 77.100 75.300 77.250 ;
        RECT 78.300 77.100 80.100 77.250 ;
        RECT 83.100 78.750 84.900 78.900 ;
        RECT 87.900 78.750 89.700 78.900 ;
        RECT 83.100 77.250 89.700 78.750 ;
        RECT 83.100 77.100 84.900 77.250 ;
        RECT 87.900 77.100 89.700 77.250 ;
        RECT 97.500 78.750 99.300 78.900 ;
        RECT 116.700 78.750 118.500 78.900 ;
        RECT 97.500 77.250 118.500 78.750 ;
        RECT 97.500 77.100 99.300 77.250 ;
        RECT 116.700 77.100 118.500 77.250 ;
        RECT 56.700 72.750 58.500 72.900 ;
        RECT 83.100 72.750 84.900 72.900 ;
        RECT 56.700 71.250 84.900 72.750 ;
        RECT 56.700 71.100 58.500 71.250 ;
        RECT 83.100 71.100 84.900 71.250 ;
        RECT 102.300 72.750 104.100 72.900 ;
        RECT 123.900 72.750 125.700 72.900 ;
        RECT 102.300 71.250 125.700 72.750 ;
        RECT 102.300 71.100 104.100 71.250 ;
        RECT 123.900 71.100 125.700 71.250 ;
        RECT 54.300 66.750 56.100 66.900 ;
        RECT 63.900 66.750 65.700 66.900 ;
        RECT 119.100 66.750 120.900 66.900 ;
        RECT 54.300 65.250 120.900 66.750 ;
        RECT 54.300 65.100 56.100 65.250 ;
        RECT 63.900 65.100 65.700 65.250 ;
        RECT 119.100 65.100 120.900 65.250 ;
        RECT 11.100 60.750 12.900 60.900 ;
        RECT 68.700 60.750 70.500 60.900 ;
        RECT 11.100 59.250 70.500 60.750 ;
        RECT 11.100 59.100 12.900 59.250 ;
        RECT 68.700 59.100 70.500 59.250 ;
        RECT 75.900 60.750 77.700 60.900 ;
        RECT 83.100 60.750 84.900 60.900 ;
        RECT 75.900 59.250 84.900 60.750 ;
        RECT 75.900 59.100 77.700 59.250 ;
        RECT 83.100 59.100 84.900 59.250 ;
        RECT 37.500 54.750 39.300 54.900 ;
        RECT 78.300 54.750 80.100 54.900 ;
        RECT 90.300 54.750 92.100 54.900 ;
        RECT 37.500 53.250 92.100 54.750 ;
        RECT 37.500 53.100 39.300 53.250 ;
        RECT 78.300 53.100 80.100 53.250 ;
        RECT 90.300 53.100 92.100 53.250 ;
        RECT 116.700 54.750 118.500 54.900 ;
        RECT 126.300 54.750 128.100 54.900 ;
        RECT 116.700 53.250 128.100 54.750 ;
        RECT 116.700 53.100 118.500 53.250 ;
        RECT 126.300 53.100 128.100 53.250 ;
        RECT 27.900 48.750 29.700 48.900 ;
        RECT 32.700 48.750 34.500 48.900 ;
        RECT 39.900 48.750 41.700 48.900 ;
        RECT 27.900 47.250 41.700 48.750 ;
        RECT 27.900 47.100 29.700 47.250 ;
        RECT 32.700 47.100 34.500 47.250 ;
        RECT 39.900 47.100 41.700 47.250 ;
        RECT 66.300 48.750 68.100 48.900 ;
        RECT 73.500 48.750 75.300 48.900 ;
        RECT 66.300 47.250 75.300 48.750 ;
        RECT 66.300 47.100 68.100 47.250 ;
        RECT 73.500 47.100 75.300 47.250 ;
        RECT 30.300 36.750 32.100 36.900 ;
        RECT 39.900 36.750 41.700 36.900 ;
        RECT 30.300 35.250 41.700 36.750 ;
        RECT 30.300 35.100 32.100 35.250 ;
        RECT 39.900 35.100 41.700 35.250 ;
        RECT 90.300 36.750 92.100 36.900 ;
        RECT 99.900 36.750 101.700 36.900 ;
        RECT 90.300 35.250 101.700 36.750 ;
        RECT 90.300 35.100 92.100 35.250 ;
        RECT 99.900 35.100 101.700 35.250 ;
        RECT 42.300 30.750 44.100 30.900 ;
        RECT 56.700 30.750 58.500 30.900 ;
        RECT 42.300 29.250 58.500 30.750 ;
        RECT 42.300 29.100 44.100 29.250 ;
        RECT 56.700 29.100 58.500 29.250 ;
        RECT 61.500 30.750 63.300 30.900 ;
        RECT 92.700 30.750 94.500 30.900 ;
        RECT 61.500 29.250 94.500 30.750 ;
        RECT 61.500 29.100 63.300 29.250 ;
        RECT 92.700 29.100 94.500 29.250 ;
        RECT 68.700 24.750 70.500 24.900 ;
        RECT 83.100 24.750 84.900 24.900 ;
        RECT 97.500 24.750 99.300 24.900 ;
        RECT 68.700 23.250 99.300 24.750 ;
        RECT 68.700 23.100 70.500 23.250 ;
        RECT 83.100 23.100 84.900 23.250 ;
        RECT 97.500 23.100 99.300 23.250 ;
        RECT 11.100 18.750 12.900 18.900 ;
        RECT 23.100 18.750 24.900 18.900 ;
        RECT 11.100 17.250 24.900 18.750 ;
        RECT 11.100 17.100 12.900 17.250 ;
        RECT 23.100 17.100 24.900 17.250 ;
        RECT 47.100 18.750 48.900 18.900 ;
        RECT 71.100 18.750 72.900 18.900 ;
        RECT 85.500 18.750 87.300 18.900 ;
        RECT 90.300 18.750 92.100 18.900 ;
        RECT 47.100 17.250 92.100 18.750 ;
        RECT 47.100 17.100 48.900 17.250 ;
        RECT 71.100 17.100 72.900 17.250 ;
        RECT 85.500 17.100 87.300 17.250 ;
        RECT 90.300 17.100 92.100 17.250 ;
        RECT 95.100 18.750 96.900 18.900 ;
        RECT 102.300 18.750 104.100 18.900 ;
        RECT 95.100 17.250 104.100 18.750 ;
        RECT 95.100 17.100 96.900 17.250 ;
        RECT 102.300 17.100 104.100 17.250 ;
        RECT 80.700 12.750 82.500 12.900 ;
        RECT 85.500 12.750 87.300 12.900 ;
        RECT 80.700 11.250 87.300 12.750 ;
        RECT 80.700 11.100 82.500 11.250 ;
        RECT 85.500 11.100 87.300 11.250 ;
        RECT 97.500 12.750 99.300 12.900 ;
        RECT 116.700 12.750 118.500 12.900 ;
        RECT 97.500 11.250 118.500 12.750 ;
        RECT 97.500 11.100 99.300 11.250 ;
        RECT 116.700 11.100 118.500 11.250 ;
  END
END processor_9_bits
END LIBRARY

